-------------------------------------------------------------------------------
-- Title      : 
-------------------------------------------------------------------------------
-- File       : PgpCardG3_DmaLoopback.vhd
-- Author     : Larry Ruckman  <ruckman@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2014-03-28
-- Last update: 2014-06-23
-- Platform   : Vivado 2013.3
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2014 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use work.StdRtlPkg.all;

-------------------------------------------------------------------------------
-- Select the PGP configuration package here
-------------------------------------------------------------------------------
use work.Pgp1p250GbpsPkg.all;

entity PgpCardG3_DmaLoopback is
   port (
      -- FLASH Interface 
      flashAddr : out   slv(25 downto 0);
      flashData : inout slv(15 downto 0);
      flashAdv  : out   sl;
      flashCe   : out   sl;
      flashOe   : out   sl;
      flashWe   : out   sl;
      -- System Signals
      sysClk     : in  sl;       -- 50 MHz
      led        : out slv(7 downto 0);
      tieToGnd   : out   slv(3 downto 0);
      tieToVdd   : out   slv(0 downto 0);
      -- PCIe Ports
      pciRstL    : in    sl;
      pciRefClkP : in    sl;            -- 100 MHz
      pciRefClkN : in    sl;            -- 100 MHz
      pciRxP     : in    slv(3 downto 0);
      pciRxN     : in    slv(3 downto 0);
      pciTxP     : out   slv(3 downto 0);
      pciTxN     : out   slv(3 downto 0));
end PgpCardG3_DmaLoopback;

architecture top_level of PgpCardG3_DmaLoopback is

begin

   PgpCardG3Core_Inst : entity work.PgpCardG3DmaLoopbackCore
      port map (
         -- FLASH Interface 
         flashAddr  => flashAddr,
         flashData  => flashData,
         flashAdv   => flashAdv,
         flashCe    => flashCe,
         flashOe    => flashOe,
         flashWe    => flashWe,
         -- System Signals
         sysClk     => sysClk,
         led        => led,
         tieToGnd   => tieToGnd,
         tieToVdd   => tieToVdd,
         -- PCIe Ports
         pciRstL    => pciRstL,
         pciRefClkP => pciRefClkP,
         pciRefClkN => pciRefClkN,
         pciRxP     => pciRxP,
         pciRxN     => pciRxN,
         pciTxP     => pciTxP,
         pciTxN     => pciTxN);   

end top_level;
